module Register(data_in, clk, en, clr, data_out);
	input [31:0] data_in;
	input clk, en, clr;
	output [31:0] data_out;
	
	My_DFFE dffe0(data_out[0],data_in[0],clk,en,clr);
	My_DFFE dffe1(data_out[1],data_in[1],clk,en,clr);
	My_DFFE dffe2(data_out[2],data_in[2],clk,en,clr);
	My_DFFE dffe3(data_out[3],data_in[3],clk,en,clr);
	My_DFFE dffe4(data_out[4],data_in[4],clk,en,clr);
	My_DFFE dffe5(data_out[5],data_in[5],clk,en,clr);
	My_DFFE dffe6(data_out[6],data_in[6],clk,en,clr);
	My_DFFE dffe7(data_out[7],data_in[7],clk,en,clr);
	My_DFFE dffe8(data_out[8],data_in[8],clk,en,clr);
	My_DFFE dffe9(data_out[9],data_in[9],clk,en,clr);
	My_DFFE dffe10(data_out[10],data_in[10],clk,en,clr);
	My_DFFE dffe11(data_out[11],data_in[11],clk,en,clr);
	My_DFFE dffe12(data_out[12],data_in[12],clk,en,clr);
	My_DFFE dffe13(data_out[13],data_in[13],clk,en,clr);
	My_DFFE dffe14(data_out[14],data_in[14],clk,en,clr);
	My_DFFE dffe15(data_out[15],data_in[15],clk,en,clr);
	My_DFFE dffe16(data_out[16],data_in[16],clk,en,clr);
	My_DFFE dffe17(data_out[17],data_in[17],clk,en,clr);
	My_DFFE dffe18(data_out[18],data_in[18],clk,en,clr);
	My_DFFE dffe19(data_out[19],data_in[19],clk,en,clr);
	My_DFFE dffe20(data_out[20],data_in[20],clk,en,clr);
	My_DFFE dffe21(data_out[21],data_in[21],clk,en,clr);
	My_DFFE dffe22(data_out[22],data_in[22],clk,en,clr);
	My_DFFE dffe23(data_out[23],data_in[23],clk,en,clr);
	My_DFFE dffe24(data_out[24],data_in[24],clk,en,clr);
	My_DFFE dffe25(data_out[25],data_in[25],clk,en,clr);
	My_DFFE dffe26(data_out[26],data_in[26],clk,en,clr);
	My_DFFE dffe27(data_out[27],data_in[27],clk,en,clr);
	My_DFFE dffe28(data_out[28],data_in[28],clk,en,clr);
	My_DFFE dffe29(data_out[29],data_in[29],clk,en,clr);
	My_DFFE dffe30(data_out[30],data_in[30],clk,en,clr);
	My_DFFE dffe31(data_out[31],data_in[31],clk,en,clr);
endmodule 