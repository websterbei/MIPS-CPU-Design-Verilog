module ThirtyTwoBitAdder(A,B,cin,S,overflow);
input [31:0] A,B;
input cin;
output [31:0] S;
output overflow;
wire cout;
wire g0,g1,g2,g3,g4,g5,g6,g7,g8,g9,g10,g11,g12,g13,g14,g15,g16,g17,g18,g19,g20,g21,g22,g23,g24,g25,g26,g27,g28,g29,g30,g31,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31;
ThirtyTwoBitCarryGenerator carryGenerator(.gm1(cin),.g0(g0),.g1(g1),.g2(g2),.g3(g3),.g4(g4),.g5(g5),.g6(g6),.g7(g7),.g8(g8),.g9(g9),.g10(g10),.g11(g11),.g12(g12),.g13(g13),.g14(g14),.g15(g15),.g16(g16),.g17(g17),.g18(g18),.g19(g19),.g20(g20),.g21(g21),.g22(g22),.g23(g23),.g24(g24),.g25(g25),.g26(g26),.g27(g27),.g28(g28),.g29(g29),.g30(g30),.g31(g31),.p0(p0),.p1(p1),.p2(p2),.p3(p3),.p4(p4),.p5(p5),.p6(p6),.p7(p7),.p8(p8),.p9(p9),.p10(p10),.p11(p11),.p12(p12),.p13(p13),.p14(p14),.p15(p15),.p16(p16),.p17(p17),.p18(p18),.p19(p19),.p20(p20),.p21(p21),.p22(p22),.p23(p23),.p24(p24),.p25(p25),.p26(p26),.p27(p27),.p28(p28),.p29(p29),.p30(p30),.p31(p31),.c1(c1),.c2(c2),.c3(c3),.c4(c4),.c5(c5),.c6(c6),.c7(c7),.c8(c8),.c9(c9),.c10(c10),.c11(c11),.c12(c12),.c13(c13),.c14(c14),.c15(c15),.c16(c16),.c17(c17),.c18(c18),.c19(c19),.c20(c20),.c21(c21),.c22(c22),.c23(c23),.c24(c24),.c25(c25),.c26(c26),.c27(c27),.c28(c28),.c29(c29),.c30(c30),.c31(c31),.c32(cout));
CarryLookaheadCell cell0(.a(A[0]), .b(B[0]), .c(cin), .s(S[0]), .g(g0), .p(p0));
CarryLookaheadCell cell1(.a(A[1]), .b(B[1]), .c(c1), .s(S[1]), .g(g1), .p(p1));
CarryLookaheadCell cell2(.a(A[2]), .b(B[2]), .c(c2), .s(S[2]), .g(g2), .p(p2));
CarryLookaheadCell cell3(.a(A[3]), .b(B[3]), .c(c3), .s(S[3]), .g(g3), .p(p3));
CarryLookaheadCell cell4(.a(A[4]), .b(B[4]), .c(c4), .s(S[4]), .g(g4), .p(p4));
CarryLookaheadCell cell5(.a(A[5]), .b(B[5]), .c(c5), .s(S[5]), .g(g5), .p(p5));
CarryLookaheadCell cell6(.a(A[6]), .b(B[6]), .c(c6), .s(S[6]), .g(g6), .p(p6));
CarryLookaheadCell cell7(.a(A[7]), .b(B[7]), .c(c7), .s(S[7]), .g(g7), .p(p7));
CarryLookaheadCell cell8(.a(A[8]), .b(B[8]), .c(c8), .s(S[8]), .g(g8), .p(p8));
CarryLookaheadCell cell9(.a(A[9]), .b(B[9]), .c(c9), .s(S[9]), .g(g9), .p(p9));
CarryLookaheadCell cell10(.a(A[10]), .b(B[10]), .c(c10), .s(S[10]), .g(g10), .p(p10));
CarryLookaheadCell cell11(.a(A[11]), .b(B[11]), .c(c11), .s(S[11]), .g(g11), .p(p11));
CarryLookaheadCell cell12(.a(A[12]), .b(B[12]), .c(c12), .s(S[12]), .g(g12), .p(p12));
CarryLookaheadCell cell13(.a(A[13]), .b(B[13]), .c(c13), .s(S[13]), .g(g13), .p(p13));
CarryLookaheadCell cell14(.a(A[14]), .b(B[14]), .c(c14), .s(S[14]), .g(g14), .p(p14));
CarryLookaheadCell cell15(.a(A[15]), .b(B[15]), .c(c15), .s(S[15]), .g(g15), .p(p15));
CarryLookaheadCell cell16(.a(A[16]), .b(B[16]), .c(c16), .s(S[16]), .g(g16), .p(p16));
CarryLookaheadCell cell17(.a(A[17]), .b(B[17]), .c(c17), .s(S[17]), .g(g17), .p(p17));
CarryLookaheadCell cell18(.a(A[18]), .b(B[18]), .c(c18), .s(S[18]), .g(g18), .p(p18));
CarryLookaheadCell cell19(.a(A[19]), .b(B[19]), .c(c19), .s(S[19]), .g(g19), .p(p19));
CarryLookaheadCell cell20(.a(A[20]), .b(B[20]), .c(c20), .s(S[20]), .g(g20), .p(p20));
CarryLookaheadCell cell21(.a(A[21]), .b(B[21]), .c(c21), .s(S[21]), .g(g21), .p(p21));
CarryLookaheadCell cell22(.a(A[22]), .b(B[22]), .c(c22), .s(S[22]), .g(g22), .p(p22));
CarryLookaheadCell cell23(.a(A[23]), .b(B[23]), .c(c23), .s(S[23]), .g(g23), .p(p23));
CarryLookaheadCell cell24(.a(A[24]), .b(B[24]), .c(c24), .s(S[24]), .g(g24), .p(p24));
CarryLookaheadCell cell25(.a(A[25]), .b(B[25]), .c(c25), .s(S[25]), .g(g25), .p(p25));
CarryLookaheadCell cell26(.a(A[26]), .b(B[26]), .c(c26), .s(S[26]), .g(g26), .p(p26));
CarryLookaheadCell cell27(.a(A[27]), .b(B[27]), .c(c27), .s(S[27]), .g(g27), .p(p27));
CarryLookaheadCell cell28(.a(A[28]), .b(B[28]), .c(c28), .s(S[28]), .g(g28), .p(p28));
CarryLookaheadCell cell29(.a(A[29]), .b(B[29]), .c(c29), .s(S[29]), .g(g29), .p(p29));
CarryLookaheadCell cell30(.a(A[30]), .b(B[30]), .c(c30), .s(S[30]), .g(g30), .p(p30));
CarryLookaheadCell cell31(.a(A[31]), .b(B[31]), .c(c31), .s(S[31]), .g(g31), .p(p31));

wire sameSign, diffSign;
xnor xnor0(sameSign, A[31], B[31]);
xor xor0(diffSign, A[31], S[31]);
and and0(overflow, sameSign, diffSign);
//xor xor0(overflow, cout, c31);
endmodule
