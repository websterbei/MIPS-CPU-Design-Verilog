module ArithmeticRightShiftByTwo(A, OUT);
input [31:0] A;
output [31:0] OUT;
assign OUT[29:0] = A[31:2];
assign OUT[31:30] = {A[31],A[31]};
endmodule 