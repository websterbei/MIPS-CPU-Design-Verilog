module ThirtyTwoBitCarryGenerator(gm1,g0,g1,g2,g3,g4,g5,g6,g7,g8,g9,g10,g11,g12,g13,g14,g15,g16,g17,g18,g19,g20,g21,g22,g23,g24,g25,g26,g27,g28,g29,g30,g31,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31,c32);
wire w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15,w16,w17,w18,w19,w20,w21,w22,w23,w24,w25,w26,w27,w28,w29,w30,w31,w32,w33,w34,w35,w36,w37,w38,w39,w40,w41,w42,w43,w44,w45,w46,w47,w48,w49,w50,w51,w52,w53,w54,w55,w56,w57,w58,w59,w60,w61,w62,w63,w64,w65,w66,w67,w68,w69,w70,w71,w72,w73,w74,w75,w76,w77,w78,w79,w80,w81,w82,w83,w84,w85,w86,w87,w88,w89,w90,w91,w92,w93,w94,w95,w96,w97,w98,w99,w100,w101,w102,w103,w104,w105,w106,w107,w108,w109,w110,w111,w112,w113,w114,w115,w116,w117,w118,w119,w120,w121,w122,w123,w124,w125,w126,w127,w128,w129,w130,w131,w132,w133,w134,w135,w136,w137,w138,w139,w140,w141,w142,w143,w144,w145,w146,w147,w148,w149,w150,w151,w152,w153,w154,w155,w156,w157,w158,w159,w160,w161,w162,w163,w164,w165,w166,w167,w168,w169,w170,w171,w172,w173,w174,w175,w176,w177,w178,w179,w180,w181,w182,w183,w184,w185,w186,w187,w188,w189,w190,w191,w192,w193,w194,w195,w196,w197,w198,w199,w200,w201,w202,w203,w204,w205,w206,w207,w208,w209,w210,w211,w212,w213,w214,w215,w216,w217,w218,w219,w220,w221,w222,w223,w224,w225,w226,w227,w228,w229,w230,w231,w232,w233,w234,w235,w236,w237,w238,w239,w240,w241,w242,w243,w244,w245,w246,w247,w248,w249,w250,w251,w252,w253,w254,w255,w256,w257,w258,w259,w260,w261,w262,w263,w264,w265,w266,w267,w268,w269,w270,w271,w272,w273,w274,w275,w276,w277,w278,w279,w280,w281,w282,w283,w284,w285,w286,w287,w288,w289,w290,w291,w292,w293,w294,w295,w296,w297,w298,w299,w300,w301,w302,w303,w304,w305,w306,w307,w308,w309,w310,w311,w312,w313,w314,w315,w316,w317,w318,w319,w320,w321,w322,w323,w324,w325,w326,w327,w328,w329,w330,w331,w332,w333,w334,w335,w336,w337,w338,w339,w340,w341,w342,w343,w344,w345,w346,w347,w348,w349,w350,w351,w352,w353,w354,w355,w356,w357,w358,w359,w360,w361,w362,w363,w364,w365,w366,w367,w368,w369,w370,w371,w372,w373,w374,w375,w376,w377,w378,w379,w380,w381,w382,w383,w384,w385,w386,w387,w388,w389,w390,w391,w392,w393,w394,w395,w396,w397,w398,w399,w400,w401,w402,w403,w404,w405,w406,w407,w408,w409,w410,w411,w412,w413,w414,w415,w416,w417,w418,w419,w420,w421,w422,w423,w424,w425,w426,w427,w428,w429,w430,w431,w432,w433,w434,w435,w436,w437,w438,w439,w440,w441,w442,w443,w444,w445,w446,w447,w448,w449,w450,w451,w452,w453,w454,w455,w456,w457,w458,w459,w460,w461,w462,w463,w464,w465,w466,w467,w468,w469,w470,w471,w472,w473,w474,w475,w476,w477,w478,w479,w480,w481,w482,w483,w484,w485,w486,w487,w488,w489,w490,w491,w492,w493,w494,w495,w496,w497,w498,w499,w500,w501,w502,w503,w504,w505,w506,w507,w508,w509,w510,w511,w512,w513,w514,w515,w516,w517,w518,w519,w520,w521,w522,w523,w524,w525,w526,w527;
input p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,gm1,g0,g1,g2,g3,g4,g5,g6,g7,g8,g9,g10,g11,g12,g13,g14,g15,g16,g17,g18,g19,g20,g21,g22,g23,g24,g25,g26,g27,g28,g29,g30,g31;
output c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31,c32;
and and0(w0,gm1,p0);
or or0(c1,g0,w0);
and and1(w1,g0,p1);
and and2(w2,gm1,p0,p1);
or or1(c2,g1,w1,w2);
and and3(w3,g1,p2);
and and4(w4,g0,p1,p2);
and and5(w5,gm1,p0,p1,p2);
or or2(c3,g2,w3,w4,w5);
and and6(w6,g2,p3);
and and7(w7,g1,p2,p3);
and and8(w8,g0,p1,p2,p3);
and and9(w9,gm1,p0,p1,p2,p3);
or or3(c4,g3,w6,w7,w8,w9);
and and10(w10,g3,p4);
and and11(w11,g2,p3,p4);
and and12(w12,g1,p2,p3,p4);
and and13(w13,g0,p1,p2,p3,p4);
and and14(w14,gm1,p0,p1,p2,p3,p4);
or or4(c5,g4,w10,w11,w12,w13,w14);
and and15(w15,g4,p5);
and and16(w16,g3,p4,p5);
and and17(w17,g2,p3,p4,p5);
and and18(w18,g1,p2,p3,p4,p5);
and and19(w19,g0,p1,p2,p3,p4,p5);
and and20(w20,gm1,p0,p1,p2,p3,p4,p5);
or or5(c6,g5,w15,w16,w17,w18,w19,w20);
and and21(w21,g5,p6);
and and22(w22,g4,p5,p6);
and and23(w23,g3,p4,p5,p6);
and and24(w24,g2,p3,p4,p5,p6);
and and25(w25,g1,p2,p3,p4,p5,p6);
and and26(w26,g0,p1,p2,p3,p4,p5,p6);
and and27(w27,gm1,p0,p1,p2,p3,p4,p5,p6);
or or6(c7,g6,w21,w22,w23,w24,w25,w26,w27);
and and28(w28,g6,p7);
and and29(w29,g5,p6,p7);
and and30(w30,g4,p5,p6,p7);
and and31(w31,g3,p4,p5,p6,p7);
and and32(w32,g2,p3,p4,p5,p6,p7);
and and33(w33,g1,p2,p3,p4,p5,p6,p7);
and and34(w34,g0,p1,p2,p3,p4,p5,p6,p7);
and and35(w35,gm1,p0,p1,p2,p3,p4,p5,p6,p7);
or or7(c8,g7,w28,w29,w30,w31,w32,w33,w34,w35);
and and36(w36,g7,p8);
and and37(w37,g6,p7,p8);
and and38(w38,g5,p6,p7,p8);
and and39(w39,g4,p5,p6,p7,p8);
and and40(w40,g3,p4,p5,p6,p7,p8);
and and41(w41,g2,p3,p4,p5,p6,p7,p8);
and and42(w42,g1,p2,p3,p4,p5,p6,p7,p8);
and and43(w43,g0,p1,p2,p3,p4,p5,p6,p7,p8);
and and44(w44,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8);
or or8(c9,g8,w36,w37,w38,w39,w40,w41,w42,w43,w44);
and and45(w45,g8,p9);
and and46(w46,g7,p8,p9);
and and47(w47,g6,p7,p8,p9);
and and48(w48,g5,p6,p7,p8,p9);
and and49(w49,g4,p5,p6,p7,p8,p9);
and and50(w50,g3,p4,p5,p6,p7,p8,p9);
and and51(w51,g2,p3,p4,p5,p6,p7,p8,p9);
and and52(w52,g1,p2,p3,p4,p5,p6,p7,p8,p9);
and and53(w53,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9);
and and54(w54,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9);
or or9(c10,g9,w45,w46,w47,w48,w49,w50,w51,w52,w53,w54);
and and55(w55,g9,p10);
and and56(w56,g8,p9,p10);
and and57(w57,g7,p8,p9,p10);
and and58(w58,g6,p7,p8,p9,p10);
and and59(w59,g5,p6,p7,p8,p9,p10);
and and60(w60,g4,p5,p6,p7,p8,p9,p10);
and and61(w61,g3,p4,p5,p6,p7,p8,p9,p10);
and and62(w62,g2,p3,p4,p5,p6,p7,p8,p9,p10);
and and63(w63,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10);
and and64(w64,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10);
and and65(w65,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10);
or or10(c11,g10,w55,w56,w57,w58,w59,w60,w61,w62,w63,w64,w65);
and and66(w66,g10,p11);
and and67(w67,g9,p10,p11);
and and68(w68,g8,p9,p10,p11);
and and69(w69,g7,p8,p9,p10,p11);
and and70(w70,g6,p7,p8,p9,p10,p11);
and and71(w71,g5,p6,p7,p8,p9,p10,p11);
and and72(w72,g4,p5,p6,p7,p8,p9,p10,p11);
and and73(w73,g3,p4,p5,p6,p7,p8,p9,p10,p11);
and and74(w74,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11);
and and75(w75,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11);
and and76(w76,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11);
and and77(w77,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11);
or or11(c12,g11,w66,w67,w68,w69,w70,w71,w72,w73,w74,w75,w76,w77);
and and78(w78,g11,p12);
and and79(w79,g10,p11,p12);
and and80(w80,g9,p10,p11,p12);
and and81(w81,g8,p9,p10,p11,p12);
and and82(w82,g7,p8,p9,p10,p11,p12);
and and83(w83,g6,p7,p8,p9,p10,p11,p12);
and and84(w84,g5,p6,p7,p8,p9,p10,p11,p12);
and and85(w85,g4,p5,p6,p7,p8,p9,p10,p11,p12);
and and86(w86,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12);
and and87(w87,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12);
and and88(w88,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12);
and and89(w89,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12);
and and90(w90,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12);
or or12(c13,g12,w78,w79,w80,w81,w82,w83,w84,w85,w86,w87,w88,w89,w90);
and and91(w91,g12,p13);
and and92(w92,g11,p12,p13);
and and93(w93,g10,p11,p12,p13);
and and94(w94,g9,p10,p11,p12,p13);
and and95(w95,g8,p9,p10,p11,p12,p13);
and and96(w96,g7,p8,p9,p10,p11,p12,p13);
and and97(w97,g6,p7,p8,p9,p10,p11,p12,p13);
and and98(w98,g5,p6,p7,p8,p9,p10,p11,p12,p13);
and and99(w99,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13);
and and100(w100,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13);
and and101(w101,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13);
and and102(w102,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13);
and and103(w103,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13);
and and104(w104,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13);
or or13(c14,g13,w91,w92,w93,w94,w95,w96,w97,w98,w99,w100,w101,w102,w103,w104);
and and105(w105,g13,p14);
and and106(w106,g12,p13,p14);
and and107(w107,g11,p12,p13,p14);
and and108(w108,g10,p11,p12,p13,p14);
and and109(w109,g9,p10,p11,p12,p13,p14);
and and110(w110,g8,p9,p10,p11,p12,p13,p14);
and and111(w111,g7,p8,p9,p10,p11,p12,p13,p14);
and and112(w112,g6,p7,p8,p9,p10,p11,p12,p13,p14);
and and113(w113,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14);
and and114(w114,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14);
and and115(w115,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14);
and and116(w116,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14);
and and117(w117,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14);
and and118(w118,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14);
and and119(w119,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14);
or or14(c15,g14,w105,w106,w107,w108,w109,w110,w111,w112,w113,w114,w115,w116,w117,w118,w119);
and and120(w120,g14,p15);
and and121(w121,g13,p14,p15);
and and122(w122,g12,p13,p14,p15);
and and123(w123,g11,p12,p13,p14,p15);
and and124(w124,g10,p11,p12,p13,p14,p15);
and and125(w125,g9,p10,p11,p12,p13,p14,p15);
and and126(w126,g8,p9,p10,p11,p12,p13,p14,p15);
and and127(w127,g7,p8,p9,p10,p11,p12,p13,p14,p15);
and and128(w128,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
and and129(w129,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
and and130(w130,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
and and131(w131,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
and and132(w132,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
and and133(w133,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
and and134(w134,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
and and135(w135,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15);
or or15(c16,g15,w120,w121,w122,w123,w124,w125,w126,w127,w128,w129,w130,w131,w132,w133,w134,w135);
and and136(w136,g15,p16);
and and137(w137,g14,p15,p16);
and and138(w138,g13,p14,p15,p16);
and and139(w139,g12,p13,p14,p15,p16);
and and140(w140,g11,p12,p13,p14,p15,p16);
and and141(w141,g10,p11,p12,p13,p14,p15,p16);
and and142(w142,g9,p10,p11,p12,p13,p14,p15,p16);
and and143(w143,g8,p9,p10,p11,p12,p13,p14,p15,p16);
and and144(w144,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and145(w145,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and146(w146,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and147(w147,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and148(w148,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and149(w149,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and150(w150,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and151(w151,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
and and152(w152,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16);
or or16(c17,g16,w136,w137,w138,w139,w140,w141,w142,w143,w144,w145,w146,w147,w148,w149,w150,w151,w152);
and and153(w153,g16,p17);
and and154(w154,g15,p16,p17);
and and155(w155,g14,p15,p16,p17);
and and156(w156,g13,p14,p15,p16,p17);
and and157(w157,g12,p13,p14,p15,p16,p17);
and and158(w158,g11,p12,p13,p14,p15,p16,p17);
and and159(w159,g10,p11,p12,p13,p14,p15,p16,p17);
and and160(w160,g9,p10,p11,p12,p13,p14,p15,p16,p17);
and and161(w161,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and162(w162,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and163(w163,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and164(w164,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and165(w165,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and166(w166,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and167(w167,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and168(w168,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and169(w169,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
and and170(w170,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17);
or or17(c18,g17,w153,w154,w155,w156,w157,w158,w159,w160,w161,w162,w163,w164,w165,w166,w167,w168,w169,w170);
and and171(w171,g17,p18);
and and172(w172,g16,p17,p18);
and and173(w173,g15,p16,p17,p18);
and and174(w174,g14,p15,p16,p17,p18);
and and175(w175,g13,p14,p15,p16,p17,p18);
and and176(w176,g12,p13,p14,p15,p16,p17,p18);
and and177(w177,g11,p12,p13,p14,p15,p16,p17,p18);
and and178(w178,g10,p11,p12,p13,p14,p15,p16,p17,p18);
and and179(w179,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and180(w180,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and181(w181,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and182(w182,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and183(w183,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and184(w184,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and185(w185,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and186(w186,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and187(w187,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and188(w188,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
and and189(w189,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18);
or or18(c19,g18,w171,w172,w173,w174,w175,w176,w177,w178,w179,w180,w181,w182,w183,w184,w185,w186,w187,w188,w189);
and and190(w190,g18,p19);
and and191(w191,g17,p18,p19);
and and192(w192,g16,p17,p18,p19);
and and193(w193,g15,p16,p17,p18,p19);
and and194(w194,g14,p15,p16,p17,p18,p19);
and and195(w195,g13,p14,p15,p16,p17,p18,p19);
and and196(w196,g12,p13,p14,p15,p16,p17,p18,p19);
and and197(w197,g11,p12,p13,p14,p15,p16,p17,p18,p19);
and and198(w198,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and199(w199,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and200(w200,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and201(w201,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and202(w202,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and203(w203,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and204(w204,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and205(w205,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and206(w206,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and207(w207,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and208(w208,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
and and209(w209,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19);
or or19(c20,g19,w190,w191,w192,w193,w194,w195,w196,w197,w198,w199,w200,w201,w202,w203,w204,w205,w206,w207,w208,w209);
and and210(w210,g19,p20);
and and211(w211,g18,p19,p20);
and and212(w212,g17,p18,p19,p20);
and and213(w213,g16,p17,p18,p19,p20);
and and214(w214,g15,p16,p17,p18,p19,p20);
and and215(w215,g14,p15,p16,p17,p18,p19,p20);
and and216(w216,g13,p14,p15,p16,p17,p18,p19,p20);
and and217(w217,g12,p13,p14,p15,p16,p17,p18,p19,p20);
and and218(w218,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and219(w219,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and220(w220,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and221(w221,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and222(w222,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and223(w223,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and224(w224,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and225(w225,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and226(w226,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and227(w227,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and228(w228,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and229(w229,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
and and230(w230,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20);
or or20(c21,g20,w210,w211,w212,w213,w214,w215,w216,w217,w218,w219,w220,w221,w222,w223,w224,w225,w226,w227,w228,w229,w230);
and and231(w231,g20,p21);
and and232(w232,g19,p20,p21);
and and233(w233,g18,p19,p20,p21);
and and234(w234,g17,p18,p19,p20,p21);
and and235(w235,g16,p17,p18,p19,p20,p21);
and and236(w236,g15,p16,p17,p18,p19,p20,p21);
and and237(w237,g14,p15,p16,p17,p18,p19,p20,p21);
and and238(w238,g13,p14,p15,p16,p17,p18,p19,p20,p21);
and and239(w239,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and240(w240,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and241(w241,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and242(w242,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and243(w243,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and244(w244,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and245(w245,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and246(w246,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and247(w247,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and248(w248,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and249(w249,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and250(w250,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and251(w251,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
and and252(w252,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21);
or or21(c22,g21,w231,w232,w233,w234,w235,w236,w237,w238,w239,w240,w241,w242,w243,w244,w245,w246,w247,w248,w249,w250,w251,w252);
and and253(w253,g21,p22);
and and254(w254,g20,p21,p22);
and and255(w255,g19,p20,p21,p22);
and and256(w256,g18,p19,p20,p21,p22);
and and257(w257,g17,p18,p19,p20,p21,p22);
and and258(w258,g16,p17,p18,p19,p20,p21,p22);
and and259(w259,g15,p16,p17,p18,p19,p20,p21,p22);
and and260(w260,g14,p15,p16,p17,p18,p19,p20,p21,p22);
and and261(w261,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and262(w262,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and263(w263,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and264(w264,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and265(w265,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and266(w266,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and267(w267,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and268(w268,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and269(w269,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and270(w270,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and271(w271,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and272(w272,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and273(w273,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and274(w274,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
and and275(w275,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22);
or or22(c23,g22,w253,w254,w255,w256,w257,w258,w259,w260,w261,w262,w263,w264,w265,w266,w267,w268,w269,w270,w271,w272,w273,w274,w275);
and and276(w276,g22,p23);
and and277(w277,g21,p22,p23);
and and278(w278,g20,p21,p22,p23);
and and279(w279,g19,p20,p21,p22,p23);
and and280(w280,g18,p19,p20,p21,p22,p23);
and and281(w281,g17,p18,p19,p20,p21,p22,p23);
and and282(w282,g16,p17,p18,p19,p20,p21,p22,p23);
and and283(w283,g15,p16,p17,p18,p19,p20,p21,p22,p23);
and and284(w284,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and285(w285,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and286(w286,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and287(w287,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and288(w288,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and289(w289,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and290(w290,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and291(w291,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and292(w292,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and293(w293,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and294(w294,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and295(w295,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and296(w296,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and297(w297,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and298(w298,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
and and299(w299,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23);
or or23(c24,g23,w276,w277,w278,w279,w280,w281,w282,w283,w284,w285,w286,w287,w288,w289,w290,w291,w292,w293,w294,w295,w296,w297,w298,w299);
and and300(w300,g23,p24);
and and301(w301,g22,p23,p24);
and and302(w302,g21,p22,p23,p24);
and and303(w303,g20,p21,p22,p23,p24);
and and304(w304,g19,p20,p21,p22,p23,p24);
and and305(w305,g18,p19,p20,p21,p22,p23,p24);
and and306(w306,g17,p18,p19,p20,p21,p22,p23,p24);
and and307(w307,g16,p17,p18,p19,p20,p21,p22,p23,p24);
and and308(w308,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and309(w309,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and310(w310,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and311(w311,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and312(w312,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and313(w313,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and314(w314,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and315(w315,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and316(w316,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and317(w317,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and318(w318,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and319(w319,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and320(w320,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and321(w321,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and322(w322,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and323(w323,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
and and324(w324,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24);
or or24(c25,g24,w300,w301,w302,w303,w304,w305,w306,w307,w308,w309,w310,w311,w312,w313,w314,w315,w316,w317,w318,w319,w320,w321,w322,w323,w324);
and and325(w325,g24,p25);
and and326(w326,g23,p24,p25);
and and327(w327,g22,p23,p24,p25);
and and328(w328,g21,p22,p23,p24,p25);
and and329(w329,g20,p21,p22,p23,p24,p25);
and and330(w330,g19,p20,p21,p22,p23,p24,p25);
and and331(w331,g18,p19,p20,p21,p22,p23,p24,p25);
and and332(w332,g17,p18,p19,p20,p21,p22,p23,p24,p25);
and and333(w333,g16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and334(w334,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and335(w335,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and336(w336,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and337(w337,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and338(w338,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and339(w339,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and340(w340,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and341(w341,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and342(w342,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and343(w343,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and344(w344,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and345(w345,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and346(w346,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and347(w347,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and348(w348,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and349(w349,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
and and350(w350,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25);
or or25(c26,g25,w325,w326,w327,w328,w329,w330,w331,w332,w333,w334,w335,w336,w337,w338,w339,w340,w341,w342,w343,w344,w345,w346,w347,w348,w349,w350);
and and351(w351,g25,p26);
and and352(w352,g24,p25,p26);
and and353(w353,g23,p24,p25,p26);
and and354(w354,g22,p23,p24,p25,p26);
and and355(w355,g21,p22,p23,p24,p25,p26);
and and356(w356,g20,p21,p22,p23,p24,p25,p26);
and and357(w357,g19,p20,p21,p22,p23,p24,p25,p26);
and and358(w358,g18,p19,p20,p21,p22,p23,p24,p25,p26);
and and359(w359,g17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and360(w360,g16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and361(w361,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and362(w362,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and363(w363,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and364(w364,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and365(w365,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and366(w366,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and367(w367,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and368(w368,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and369(w369,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and370(w370,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and371(w371,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and372(w372,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and373(w373,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and374(w374,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and375(w375,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and376(w376,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
and and377(w377,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26);
or or26(c27,g26,w351,w352,w353,w354,w355,w356,w357,w358,w359,w360,w361,w362,w363,w364,w365,w366,w367,w368,w369,w370,w371,w372,w373,w374,w375,w376,w377);
and and378(w378,g26,p27);
and and379(w379,g25,p26,p27);
and and380(w380,g24,p25,p26,p27);
and and381(w381,g23,p24,p25,p26,p27);
and and382(w382,g22,p23,p24,p25,p26,p27);
and and383(w383,g21,p22,p23,p24,p25,p26,p27);
and and384(w384,g20,p21,p22,p23,p24,p25,p26,p27);
and and385(w385,g19,p20,p21,p22,p23,p24,p25,p26,p27);
and and386(w386,g18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and387(w387,g17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and388(w388,g16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and389(w389,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and390(w390,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and391(w391,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and392(w392,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and393(w393,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and394(w394,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and395(w395,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and396(w396,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and397(w397,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and398(w398,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and399(w399,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and400(w400,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and401(w401,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and402(w402,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and403(w403,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and404(w404,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
and and405(w405,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27);
or or27(c28,g27,w378,w379,w380,w381,w382,w383,w384,w385,w386,w387,w388,w389,w390,w391,w392,w393,w394,w395,w396,w397,w398,w399,w400,w401,w402,w403,w404,w405);
and and406(w406,g27,p28);
and and407(w407,g26,p27,p28);
and and408(w408,g25,p26,p27,p28);
and and409(w409,g24,p25,p26,p27,p28);
and and410(w410,g23,p24,p25,p26,p27,p28);
and and411(w411,g22,p23,p24,p25,p26,p27,p28);
and and412(w412,g21,p22,p23,p24,p25,p26,p27,p28);
and and413(w413,g20,p21,p22,p23,p24,p25,p26,p27,p28);
and and414(w414,g19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and415(w415,g18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and416(w416,g17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and417(w417,g16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and418(w418,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and419(w419,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and420(w420,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and421(w421,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and422(w422,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and423(w423,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and424(w424,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and425(w425,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and426(w426,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and427(w427,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and428(w428,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and429(w429,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and430(w430,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and431(w431,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and432(w432,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and433(w433,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
and and434(w434,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28);
or or28(c29,g28,w406,w407,w408,w409,w410,w411,w412,w413,w414,w415,w416,w417,w418,w419,w420,w421,w422,w423,w424,w425,w426,w427,w428,w429,w430,w431,w432,w433,w434);
and and435(w435,g28,p29);
and and436(w436,g27,p28,p29);
and and437(w437,g26,p27,p28,p29);
and and438(w438,g25,p26,p27,p28,p29);
and and439(w439,g24,p25,p26,p27,p28,p29);
and and440(w440,g23,p24,p25,p26,p27,p28,p29);
and and441(w441,g22,p23,p24,p25,p26,p27,p28,p29);
and and442(w442,g21,p22,p23,p24,p25,p26,p27,p28,p29);
and and443(w443,g20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and444(w444,g19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and445(w445,g18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and446(w446,g17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and447(w447,g16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and448(w448,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and449(w449,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and450(w450,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and451(w451,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and452(w452,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and453(w453,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and454(w454,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and455(w455,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and456(w456,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and457(w457,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and458(w458,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and459(w459,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and460(w460,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and461(w461,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and462(w462,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and463(w463,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
and and464(w464,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29);
or or29(c30,g29,w435,w436,w437,w438,w439,w440,w441,w442,w443,w444,w445,w446,w447,w448,w449,w450,w451,w452,w453,w454,w455,w456,w457,w458,w459,w460,w461,w462,w463,w464);
and and465(w465,g29,p30);
and and466(w466,g28,p29,p30);
and and467(w467,g27,p28,p29,p30);
and and468(w468,g26,p27,p28,p29,p30);
and and469(w469,g25,p26,p27,p28,p29,p30);
and and470(w470,g24,p25,p26,p27,p28,p29,p30);
and and471(w471,g23,p24,p25,p26,p27,p28,p29,p30);
and and472(w472,g22,p23,p24,p25,p26,p27,p28,p29,p30);
and and473(w473,g21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and474(w474,g20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and475(w475,g19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and476(w476,g18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and477(w477,g17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and478(w478,g16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and479(w479,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and480(w480,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and481(w481,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and482(w482,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and483(w483,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and484(w484,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and485(w485,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and486(w486,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and487(w487,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and488(w488,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and489(w489,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and490(w490,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and491(w491,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and492(w492,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and493(w493,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and494(w494,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
and and495(w495,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30);
or or30(c31,g30,w465,w466,w467,w468,w469,w470,w471,w472,w473,w474,w475,w476,w477,w478,w479,w480,w481,w482,w483,w484,w485,w486,w487,w488,w489,w490,w491,w492,w493,w494,w495);
and and496(w496,g30,p31);
and and497(w497,g29,p30,p31);
and and498(w498,g28,p29,p30,p31);
and and499(w499,g27,p28,p29,p30,p31);
and and500(w500,g26,p27,p28,p29,p30,p31);
and and501(w501,g25,p26,p27,p28,p29,p30,p31);
and and502(w502,g24,p25,p26,p27,p28,p29,p30,p31);
and and503(w503,g23,p24,p25,p26,p27,p28,p29,p30,p31);
and and504(w504,g22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and505(w505,g21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and506(w506,g20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and507(w507,g19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and508(w508,g18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and509(w509,g17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and510(w510,g16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and511(w511,g15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and512(w512,g14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and513(w513,g13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and514(w514,g12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and515(w515,g11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and516(w516,g10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and517(w517,g9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and518(w518,g8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and519(w519,g7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and520(w520,g6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and521(w521,g5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and522(w522,g4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and523(w523,g3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and524(w524,g2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and525(w525,g1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and526(w526,g0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
and and527(w527,gm1,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31);
or or31(c32,g31,w496,w497,w498,w499,w500,w501,w502,w503,w504,w505,w506,w507,w508,w509,w510,w511,w512,w513,w514,w515,w516,w517,w518,w519,w520,w521,w522,w523,w524,w525,w526,w527);
endmodule
